LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.MATH_REAL.LOG2;
USE IEEE.MATH_REAL.CEIL;

--THIS VERSION USES TWO POINTER AND WRITING AND READING SIMULTANEOUSLY
ENTITY KASO_BUFF IS
GENERIC(
			K: INTEGER:=4; 
			N: INTEGER :=10; 
			PIXEL:INTEGER:=30
			);
PORT(
	  SAMPLE					: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	  READY					: IN STD_LOGIC;
	  CLK,RESET				: IN STD_LOGIC;
	  ENERGY					: OUT STD_LOGIC_VECTOR(2*N-1 DOWNTO 0);
	  INDEXW					: IN UNSIGNED(INTEGER(CEIL(LOG2(REAL((K*PIXEL+1)))))-1 DOWNTO 0);
	  INDEXK					: IN UNSIGNED(INTEGER(CEIL(LOG2(REAL((K*PIXEL+1)))))-1 DOWNTO 0)
	 
	  );
END ENTITY KASO_BUFF;

ARCHITECTURE RTL OF KASO_BUFF IS
TYPE MAT IS ARRAY(0 TO K*PIXEL) OF STD_LOGIC_VECTOR(N-1 DOWNTO 0);
SIGNAL Q													: MAT;
SIGNAL SQ												: SIGNED (2*N-1 DOWNTO 0);
SIGNAL MK												: SIGNED	(N-1 DOWNTO 0);





BEGIN




MEMORY:PROCESS(CLK,RESET) 
BEGIN
IF(RESET='0') THEN
	Q<=(OTHERS=>(OTHERS=>'0'));
ELSIF(RISING_EDGE(CLK)) THEN
 
 	Q(TO_INTEGER(INDEXW))<=SAMPLE;
	
END IF;

END PROCESS MEMORY;




  
 MK<=SIGNED(Q(TO_INTEGER(INDEXK)))-SIGNED(Q(TO_INTEGER(INDEXW))); --X(N)-X(N-K)
 SQ<=SIGNED(Q(TO_INTEGER(INDEXK)))*MK; --X(N) (X(N)-X(N-K))
 ENERGY<=STD_LOGIC_VECTOR(SQ(2*N-1 DOWNTO 0)) WHEN (READY='0') ELSE (OTHERS=>'0');

	
END ARCHITECTURE RTL;
