LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.MATH_REAL.LOG2;
USE IEEE.MATH_REAL.CEIL;

USE WORK.VHDLTOOL.ALL;

--BUFFERIZED R/W SIMULTANEOUS
ENTITY SMOOTHING_BUFF IS
GENERIC(
			CHANNEL	: INTEGER:=30; 
			K			: INTEGER:=4; 
			N			: INTEGER:=10
			);
PORT( 
		SAMPLE				: IN STD_LOGIC_VECTOR(2*N-1 DOWNTO 0); --Q19.0
		CLK,RESET			: IN STD_LOGIC;
		INDEXR				: IN POINTERS (0 TO 4*K);
		INDEXW				: IN UNSIGNED(INTEGER(CEIL(LOG2(REAL(4*K*CHANNEL+1))))-1 DOWNTO 0);
		READY					: IN STD_LOGIC;
		SMOOTHED				: OUT STD_LOGIC_VECTOR(2*N-1 DOWNTO 0) --Q19.0
		);
END SMOOTHING_BUFF;

ARCHITECTURE RTL OF SMOOTHING_BUFF IS 
-- HAMMING FIR COEFFICIENT L=64, K=4 Q9.0
CONSTANT B0: SIGNED (N-1 DOWNTO 0) := TO_SIGNED(5,10);
CONSTANT B1: SIGNED (N-1 DOWNTO 0) := TO_SIGNED(7,10);
CONSTANT B2: SIGNED (N-1 DOWNTO 0) := TO_SIGNED(13,10);
CONSTANT B3: SIGNED (N-1 DOWNTO 0) := TO_SIGNED(21,10);
CONSTANT B4: SIGNED (N-1 DOWNTO 0) := TO_SIGNED(32,10);
CONSTANT B5: SIGNED (N-1 DOWNTO 0) := TO_SIGNED(42,10);
CONSTANT B6: SIGNED (N-1 DOWNTO 0) := TO_SIGNED(51,10);
CONSTANT B7: SIGNED (N-1 DOWNTO 0) := TO_SIGNED(57,10);
CONSTANT B8: SIGNED (N-1 DOWNTO 0) := TO_SIGNED(59,10);




TYPE MAT IS ARRAY (0 TO 4*K*CHANNEL) OF STD_LOGIC_VECTOR(2*N-1 DOWNTO 0);
SIGNAL Q: MAT;

BEGIN


--DEALY BLOCK
DELAYBLOCK:PROCESS(CLK,RESET)
BEGIN
IF (RESET='0') THEN
	Q<=(OTHERS=>(OTHERS=>'0'));
ELSIF (RISING_EDGE(CLK)) THEN
		Q(TO_INTEGER(INDEXW))<=SAMPLE;
END IF;

END PROCESS DELAYBLOCK;

PROCESS(INDEXR,Q,READY)
VARIABLE SUM,M1,M2,M3,M4,M5,M6,M7,M8,M9,M10,M11,M12,M13,M14,M15,M16,M17: SIGNED(3*N-1 DOWNTO 0) ; --Q29.0

BEGIN
-- MULTIPLICATIONS
IF(READY='0') THEN
	M1:=SIGNED(Q(TO_INTEGER(INDEXR(16))))*B0;
	M2:=SIGNED(Q(TO_INTEGER(INDEXR(15))))*B1;
	M3:=SIGNED(Q(TO_INTEGER(INDEXR(14))))*B2;
	M4:=SIGNED(Q(TO_INTEGER(INDEXR(13))))*B3;
	M5:=SIGNED(Q(TO_INTEGER(INDEXR(12))))*B4;
	M6:=SIGNED(Q(TO_INTEGER(INDEXR(11))))*B5;
	M7:=SIGNED(Q(TO_INTEGER(INDEXR(10))))*B6;
	M8:=SIGNED(Q(TO_INTEGER(INDEXR(9))))*B7;
	M9:=SIGNED(Q(TO_INTEGER(INDEXR(8))))*B8;
	M10:=SIGNED(Q(TO_INTEGER(INDEXR(7))))*B7;
	M11:=SIGNED(Q(TO_INTEGER(INDEXR(6))))*B6;
	M12:=SIGNED(Q(TO_INTEGER(INDEXR(5))))*B5;
	M13:=SIGNED(Q(TO_INTEGER(INDEXR(4))))*B4;
	M14:=SIGNED(Q(TO_INTEGER(INDEXR(3))))*B3;
	M15:=SIGNED(Q(TO_INTEGER(INDEXR(2))))*B2;
	M16:=SIGNED(Q(TO_INTEGER(INDEXR(1))))*B1;
	M17:=SIGNED(Q(TO_INTEGER(INDEXR(0))))*B0;
	
	
	SUM:= M1+M2+M3+M4+M5+M6+M7+M8+M9+M10+M11+M12+M13+M14+M15+M16+M17;
	SMOOTHED<=STD_LOGIC_VECTOR(SUM(3*N-2 DOWNTO N-1)); --Q19.0
ELSE
	SMOOTHED<=(OTHERS=>'0'); --Q19.0
END IF;
END PROCESS;




END ARCHITECTURE RTL;
