LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.MATH_REAL.LOG2;
USE IEEE.MATH_REAL.CEIL;

--VERSION 2 USED TO RECOVER CLOCK STROKES WRITING AND READING IN SIMULATANEA DELLA STESSA LOCAZIONE ATTENZIONE
ENTITY KASO_CONTROLLER IS
GENERIC (
			K       : INTEGER:=4; 
			PIXEL	: INTEGER
			);
PORT 	(	
			CLK,RESET,ENABLE	: IN STD_LOGIC;
			READY			: OUT STD_LOGIC;
			INDEXW			: OUT UNSIGNED(INTEGER(CEIL(LOG2(REAL(K*PIXEL+1))))-1 DOWNTO 0);
			INDEXK			: OUT UNSIGNED(INTEGER(CEIL(LOG2(REAL(K*PIXEL+1))))-1 DOWNTO 0)
);
END ENTITY KASO_CONTROLLER;

ARCHITECTURE RTL OF KASO_CONTROLLER IS
SIGNAL READY_TMP: STD_LOGIC;
BEGIN

-----POINTERS LOGIC
WRITEMEM:PROCESS(CLK,RESET) 
VARIABLE CNT_NEW: UNSIGNED( INTEGER(CEIL(LOG2(REAL(K*PIXEL+1))))-1 DOWNTO 0);
BEGIN
IF(RESET='0') THEN
	CNT_NEW:=(OTHERS=>'0');
	READY_TMP<='1';
ELSIF(RISING_EDGE(CLK)) THEN
 IF(ENABLE='0') THEN
	
	 CNT_NEW:=CNT_NEW+1;
		
	IF(CNT_NEW=K*PIXEL+1) THEN
				CNT_NEW:=(OTHERS=>'0');
				READY_TMP<='0';
			END IF;
	
	
END IF;
END IF;
INDEXW<=CNT_NEW;
END PROCESS WRITEMEM;

READY<=READY_TMP;


INDEXINGOLDSAMPLEW:PROCESS(CLK,RESET) 
VARIABLE CNT_NEW: UNSIGNED( INTEGER(CEIL(LOG2(REAL(K*PIXEL+1))))-1 DOWNTO 0);
BEGIN
IF(RESET='0') THEN
	CNT_NEW:=TO_UNSIGNED((K*PIXEL),CNT_NEW'LENGTH);
ELSIF(RISING_EDGE(CLK)) THEN
 IF(READY_TMP='0') THEN
	
	 CNT_NEW:=CNT_NEW+1;
		
	 IF(CNT_NEW=K*PIXEL+1) THEN
	 
			CNT_NEW:=(OTHERS=>'0');
				
	 END IF;
	
	
 END IF;
END IF;
INDEXK<=CNT_NEW;
END PROCESS INDEXINGOLDSAMPLEW;






END ARCHITECTURE RTL; 
