LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

--THE SCRIPT CONTAINS AT THE END THE ADDITIONAL MODULES USED INTO THE MAIN ONE.



ENTITY STATIC_MEDIAN IS 
PORT(
		SAMPLE: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		READY	: OUT STD_LOGIC;
		CLK,RESET,ENABLE: IN STD_LOGIC;
		MEDIAN: OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
		
		);
END ENTITY STATIC_MEDIAN;

ARCHITECTURE RTL OF STATIC_MEDIAN IS
-- COMPONENT INSTANCES
COMPONENT NODEBIN IS
	 GENERIC(
					MEDIAN_INDEX:INTEGER;
					MEDIAN_LEN: INTEGER
				);
	 PORT( 
				SEL: IN STD_LOGIC;
				CLK,RESET,CLEAR,ENABLE: IN STD_LOGIC;
				GTMED: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
			 );
	END COMPONENT NODEBIN;
	
COMPONENT LASTNODEBIN IS 
GENERIC(
			MEDIAN_INDEX:INTEGER:=32; 
			MEDIAN_LEN: INTEGER:=64
			);
	PORT( 
			SEL: IN STD_LOGIC;
			CLK,RESET,ENABLE:IN STD_LOGIC;
			COUT: OUT STD_LOGIC;
			GTMED: OUT STD_LOGIC_VECTOR(1 DOWNTO 0) --USING TO BIT ONE FOR 31TH INDEX AND THE LSB FOR 32TH BIT
		);
END COMPONENT LASTNODEBIN;

COMPONENT SELECTORBIN IS
	 PORT(
				SEL: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
				ENABLE:IN STD_LOGIC;
				LUT_OUT: OUT STD_LOGIC_VECTOR (511 DOWNTO 0)
			);
END COMPONENT SELECTORBIN;

COMPONENT PRIORENCMEDIAN IS 
	 PORT(
				GTMED_S: IN STD_LOGIC_VECTOR(511 DOWNTO 0);
				MEDIAN: OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
		   );
END COMPONENT PRIORENCMEDIAN;


--SIGNAL DECLARATIONS
SIGNAL DECODED: STD_LOGIC_VECTOR(511 DOWNTO 0);
TYPE INDEXM IS ARRAY (0 TO 511) OF STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL GTMED_S: INDEXM;

SIGNAL EVENINDEX,ODDINDEX: STD_LOGIC_VECTOR(511 DOWNTO 0);
SIGNAL Q,POSITIVO: STD_LOGIC_VECTOR(8 DOWNTO 0);
CONSTANT C: UNSIGNED(3 DOWNTO 0):=TO_UNSIGNED(11,4); --U-1.4 11 0.6745 TRUE VAL 0.6745
SIGNAL TMP1,TMP2,SUM: STD_LOGIC_VECTOR(8 DOWNTO 0); 
SIGNAL SUMTMP: UNSIGNED(9 DOWNTO 0);
SIGNAL CNT:STD_LOGIC;
SIGNAL MQ: UNSIGNED(Q'LENGTH+C'LENGTH-1 DOWNTO 0);
SIGNAL POS_TEMP: SIGNED(9 DOWNTO 0);

BEGIN

POS_TEMP<=ABS(SIGNED(SAMPLE));
POSITIVO<=STD_LOGIC_VECTOR(POS_TEMP(8 DOWNTO 0));


SAMPLING: PROCESS(CLK) --IT MAY BE CHANGED DEPENDING ON THE BLOCK BEFORE IT.
BEGIN
IF(RISING_EDGE(CLK)) THEN
	IF(RESET='0') THEN
		Q<=(OTHERS=>'0');
	 ELSE
		Q<=POSITIVO;
	END IF;
		
END IF;
END PROCESS SAMPLING;

DECODER: SELECTORBIN PORT MAP(SEL=>Q,ENABLE=>ENABLE,LUT_OUT=>DECODED);  --RESET USED AS ENABLE SIGNAL

BINS:FOR I IN 0 TO 511 GENERATE
	FIRSTBINS: IF I<511 GENERATE
		BINELEM: NODEBIN 	GENERIC MAP(32,64)
								PORT MAP(SEL=>DECODED(I),CLK=>CLK,RESET=>RESET,CLEAR=>CNT,ENABLE=>ENABLE,GTMED=>GTMED_S(I));
					END GENERATE FIRSTBINS;
			LAST:IF (I=511) GENERATE
			         LASTBIN: LASTNODEBIN GENERIC MAP(32,64)
									PORT MAP(SEL=>DECODED(I),CLK=>CLK,RESET=>RESET,ENABLE=>ENABLE,COUT=>CNT,GTMED=>GTMED_S(I));
					END GENERATE LAST;
		END GENERATE BINS;
		
SLICINGARRAY:PROCESS(GTMED_S)
	VARIABLE TMP1: STD_LOGIC_VECTOR(GTMED_S'REVERSE_RANGE);
	VARIABLE TMP2: STD_LOGIC_VECTOR(GTMED_S'REVERSE_RANGE);
BEGIN
	FOR I IN GTMED_S'REVERSE_RANGE LOOP
		TMP1(I):=GTMED_S(I)(1);
		TMP2(I):=GTMED_S(I)(0);
	END LOOP;
		EVENINDEX<=TMP1;
		ODDINDEX<=TMP2;
END PROCESS SLICINGARRAY;



LASTBLOCKEVENDINX: PRIORENCMEDIAN PORT MAP(GTMED_S=>EVENINDEX,MEDIAN=>TMP1);
LASTBLOCKEVODD: PRIORENCMEDIAN PORT MAP(GTMED_S=>ODDINDEX,MEDIAN=>TMP2);

SUMTMP<=('0'& UNSIGNED(TMP1))+('0'& UNSIGNED(TMP2));

MQ<=SUMTMP(SUMTMP'HIGH DOWNTO 1)*C;

SUM<=STD_LOGIC_VECTOR(MQ(MQ'LENGTH-1 DOWNTO 4));

UPDATE:PROCESS(CLK,RESET)
BEGIN
IF (RESET='0') THEN
	MEDIAN<=(OTHERS=>'0');
	READY<='1';
ELSIF(RISING_EDGE(CLK)) THEN
  IF (CNT='1') THEN
    MEDIAN<=SUM;
	 READY<='0';
  END IF;
END IF;
END PROCESS UPDATE;	
	

END ARCHITECTURE RTL;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY LASTNODEBIN IS 
GENERIC(MEDIAN_INDEX:INTEGER:=32; MEDIAN_LEN: INTEGER:=64);
PORT( SEL: IN STD_LOGIC;
		CLK,RESET,ENABLE:IN STD_LOGIC;
		COUT: OUT STD_LOGIC;
		GTMED: OUT STD_LOGIC_VECTOR(1 DOWNTO 0) --USING TO BIT ONE FOR 31TH INDEX AND THE LSB FOR 32TH BIT
		);
END ENTITY LASTNODEBIN;

ARCHITECTURE RTL OF LASTNODEBIN IS 
SIGNAL Y  : UNSIGNED(5 DOWNTO 0);
SIGNAL SUM: UNSIGNED(5 DOWNTO 0);
BEGIN

Y<=SUM+1 WHEN (SEL='1') ELSE SUM;

UPDATE: PROCESS(CLK,RESET)
VARIABLE C:STD_LOGIC;
BEGIN
IF (RESET='0') THEN
	SUM<=(OTHERS=>'0');
	C:='0';
	GTMED<=(OTHERS=>'0');

ELSIF (RISING_EDGE(CLK)) THEN
   IF(ENABLE='0') THEN  
		
		 SUM<=Y;
		 
		 IF(SUM>MEDIAN_INDEX-1) THEN
		  GTMED(1)<='1';
		  IF (SUM>MEDIAN_INDEX) THEN
		  GTMED(0)<='1';
		  IF (SUM=MEDIAN_LEN-1) THEN
		   C:='1';
			SUM<=(OTHERS=>'0');
		   END IF;
		  END IF;
		 ELSE 
		  GTMED<="00";
		  C:='0';
		END IF;
	END IF;
END IF;
COUT<=C;
END PROCESS UPDATE;
END ARCHITECTURE RTL;




LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY NODEBIN IS 
GENERIC(MEDIAN_INDEX:INTEGER:=32; MEDIAN_LEN: INTEGER:=64);
PORT( SEL: IN STD_LOGIC;
		CLK,RESET,CLEAR,ENABLE:IN STD_LOGIC;
		GTMED: OUT STD_LOGIC_VECTOR(1 DOWNTO 0) --USING TO BIT ONE FOR 31TH INDEX AND THE LSB FOR 32TH BIT
		);
END ENTITY NODEBIN;

ARCHITECTURE RTL OF NODEBIN IS 
SIGNAL Y  : UNSIGNED(5 DOWNTO 0);
SIGNAL SUM: UNSIGNED(5 DOWNTO 0);
BEGIN

Y<=SUM+1 WHEN (SEL='1') ELSE SUM;

UPDATE: PROCESS(CLK,RESET)
BEGIN
IF (RESET='0') THEN
	SUM<=(OTHERS=>'0');
	GTMED<=(OTHERS=>'0');

ELSIF (RISING_EDGE(CLK)) THEN
   IF(ENABLE='0') THEN  
		IF(CLEAR='1') THEN
			SUM<=(OTHERS=>'0');
		ELSE
		 SUM<=Y;
		 END IF;
		 IF(SUM>MEDIAN_INDEX-1) THEN
		  GTMED(1)<='1';
		  IF (SUM>MEDIAN_INDEX) THEN
		   GTMED(0)<='1';
		 END IF;
		 ELSE 
		  GTMED<="00";
		END IF;
	END IF;
END IF;
END PROCESS UPDATE;
END ARCHITECTURE RTL;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY PRIORENCMEDIAN IS 
PORT(GTMED_S: IN STD_LOGIC_VECTOR(511 DOWNTO 0);
	  MEDIAN: OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	  );
END ENTITY PRIORENCMEDIAN;

ARCHITECTURE RTL OF PRIORENCMEDIAN IS

BEGIN


	MEDIAN <= STD_LOGIC_VECTOR(TO_UNSIGNED(0,9)) WHEN GTMED_S(0)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(1,9)) WHEN GTMED_S(1)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(2,9)) WHEN GTMED_S(2)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(3,9)) WHEN GTMED_S(3)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(4,9)) WHEN GTMED_S(4)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(5,9)) WHEN GTMED_S(5)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(6,9)) WHEN GTMED_S(6)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(7,9)) WHEN GTMED_S(7)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(8,9)) WHEN GTMED_S(8)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(9,9)) WHEN GTMED_S(9)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(10,9)) WHEN GTMED_S(10)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(11,9)) WHEN GTMED_S(11)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(12,9)) WHEN GTMED_S(12)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(13,9)) WHEN GTMED_S(13)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(14,9)) WHEN GTMED_S(14)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(15,9)) WHEN GTMED_S(15)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(16,9)) WHEN GTMED_S(16)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(17,9)) WHEN GTMED_S(17)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(18,9)) WHEN GTMED_S(18)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(19,9)) WHEN GTMED_S(19)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(20,9)) WHEN GTMED_S(20)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(21,9)) WHEN GTMED_S(21)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(22,9)) WHEN GTMED_S(22)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(23,9)) WHEN GTMED_S(23)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(24,9)) WHEN GTMED_S(24)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(25,9)) WHEN GTMED_S(25)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(26,9)) WHEN GTMED_S(26)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(27,9)) WHEN GTMED_S(27)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(28,9)) WHEN GTMED_S(28)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(29,9)) WHEN GTMED_S(29)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(30,9)) WHEN GTMED_S(30)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(31,9)) WHEN GTMED_S(31)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(32,9)) WHEN GTMED_S(32)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(33,9)) WHEN GTMED_S(33)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(34,9)) WHEN GTMED_S(34)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(35,9)) WHEN GTMED_S(35)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(36,9)) WHEN GTMED_S(36)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(37,9)) WHEN GTMED_S(37)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(38,9)) WHEN GTMED_S(38)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(39,9)) WHEN GTMED_S(39)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(40,9)) WHEN GTMED_S(40)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(41,9)) WHEN GTMED_S(41)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(42,9)) WHEN GTMED_S(42)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(43,9)) WHEN GTMED_S(43)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(44,9)) WHEN GTMED_S(44)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(45,9)) WHEN GTMED_S(45)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(46,9)) WHEN GTMED_S(46)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(47,9)) WHEN GTMED_S(47)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(48,9)) WHEN GTMED_S(48)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(49,9)) WHEN GTMED_S(49)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(50,9)) WHEN GTMED_S(50)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(51,9)) WHEN GTMED_S(51)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(52,9)) WHEN GTMED_S(52)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(53,9)) WHEN GTMED_S(53)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(54,9)) WHEN GTMED_S(54)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(55,9)) WHEN GTMED_S(55)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(56,9)) WHEN GTMED_S(56)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(57,9)) WHEN GTMED_S(57)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(58,9)) WHEN GTMED_S(58)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(59,9)) WHEN GTMED_S(59)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(60,9)) WHEN GTMED_S(60)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(61,9)) WHEN GTMED_S(61)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(62,9)) WHEN GTMED_S(62)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(63,9)) WHEN GTMED_S(63)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(64,9)) WHEN GTMED_S(64)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(65,9)) WHEN GTMED_S(65)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(66,9)) WHEN GTMED_S(66)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(67,9)) WHEN GTMED_S(67)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(68,9)) WHEN GTMED_S(68)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(69,9)) WHEN GTMED_S(69)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(70,9)) WHEN GTMED_S(70)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(71,9)) WHEN GTMED_S(71)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(72,9)) WHEN GTMED_S(72)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(73,9)) WHEN GTMED_S(73)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(74,9)) WHEN GTMED_S(74)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(75,9)) WHEN GTMED_S(75)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(76,9)) WHEN GTMED_S(76)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(77,9)) WHEN GTMED_S(77)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(78,9)) WHEN GTMED_S(78)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(79,9)) WHEN GTMED_S(79)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(80,9)) WHEN GTMED_S(80)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(81,9)) WHEN GTMED_S(81)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(82,9)) WHEN GTMED_S(82)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(83,9)) WHEN GTMED_S(83)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(84,9)) WHEN GTMED_S(84)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(85,9)) WHEN GTMED_S(85)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(86,9)) WHEN GTMED_S(86)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(87,9)) WHEN GTMED_S(87)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(88,9)) WHEN GTMED_S(88)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(89,9)) WHEN GTMED_S(89)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(90,9)) WHEN GTMED_S(90)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(91,9)) WHEN GTMED_S(91)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(92,9)) WHEN GTMED_S(92)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(93,9)) WHEN GTMED_S(93)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(94,9)) WHEN GTMED_S(94)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(95,9)) WHEN GTMED_S(95)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(96,9)) WHEN GTMED_S(96)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(97,9)) WHEN GTMED_S(97)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(98,9)) WHEN GTMED_S(98)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(99,9)) WHEN GTMED_S(99)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(100,9)) WHEN GTMED_S(100)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(101,9)) WHEN GTMED_S(101)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(102,9)) WHEN GTMED_S(102)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(103,9)) WHEN GTMED_S(103)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(104,9)) WHEN GTMED_S(104)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(105,9)) WHEN GTMED_S(105)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(106,9)) WHEN GTMED_S(106)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(107,9)) WHEN GTMED_S(107)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(108,9)) WHEN GTMED_S(108)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(109,9)) WHEN GTMED_S(109)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(110,9)) WHEN GTMED_S(110)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(111,9)) WHEN GTMED_S(111)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(112,9)) WHEN GTMED_S(112)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(113,9)) WHEN GTMED_S(113)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(114,9)) WHEN GTMED_S(114)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(115,9)) WHEN GTMED_S(115)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(116,9)) WHEN GTMED_S(116)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(117,9)) WHEN GTMED_S(117)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(118,9)) WHEN GTMED_S(118)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(119,9)) WHEN GTMED_S(119)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(120,9)) WHEN GTMED_S(120)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(121,9)) WHEN GTMED_S(121)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(122,9)) WHEN GTMED_S(122)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(123,9)) WHEN GTMED_S(123)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(124,9)) WHEN GTMED_S(124)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(125,9)) WHEN GTMED_S(125)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(126,9)) WHEN GTMED_S(126)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(127,9)) WHEN GTMED_S(127)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(128,9)) WHEN GTMED_S(128)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(129,9)) WHEN GTMED_S(129)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(130,9)) WHEN GTMED_S(130)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(131,9)) WHEN GTMED_S(131)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(132,9)) WHEN GTMED_S(132)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(133,9)) WHEN GTMED_S(133)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(134,9)) WHEN GTMED_S(134)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(135,9)) WHEN GTMED_S(135)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(136,9)) WHEN GTMED_S(136)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(137,9)) WHEN GTMED_S(137)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(138,9)) WHEN GTMED_S(138)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(139,9)) WHEN GTMED_S(139)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(140,9)) WHEN GTMED_S(140)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(141,9)) WHEN GTMED_S(141)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(142,9)) WHEN GTMED_S(142)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(143,9)) WHEN GTMED_S(143)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(144,9)) WHEN GTMED_S(144)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(145,9)) WHEN GTMED_S(145)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(146,9)) WHEN GTMED_S(146)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(147,9)) WHEN GTMED_S(147)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(148,9)) WHEN GTMED_S(148)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(149,9)) WHEN GTMED_S(149)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(150,9)) WHEN GTMED_S(150)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(151,9)) WHEN GTMED_S(151)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(152,9)) WHEN GTMED_S(152)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(153,9)) WHEN GTMED_S(153)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(154,9)) WHEN GTMED_S(154)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(155,9)) WHEN GTMED_S(155)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(156,9)) WHEN GTMED_S(156)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(157,9)) WHEN GTMED_S(157)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(158,9)) WHEN GTMED_S(158)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(159,9)) WHEN GTMED_S(159)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(160,9)) WHEN GTMED_S(160)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(161,9)) WHEN GTMED_S(161)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(162,9)) WHEN GTMED_S(162)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(163,9)) WHEN GTMED_S(163)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(164,9)) WHEN GTMED_S(164)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(165,9)) WHEN GTMED_S(165)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(166,9)) WHEN GTMED_S(166)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(167,9)) WHEN GTMED_S(167)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(168,9)) WHEN GTMED_S(168)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(169,9)) WHEN GTMED_S(169)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(170,9)) WHEN GTMED_S(170)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(171,9)) WHEN GTMED_S(171)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(172,9)) WHEN GTMED_S(172)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(173,9)) WHEN GTMED_S(173)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(174,9)) WHEN GTMED_S(174)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(175,9)) WHEN GTMED_S(175)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(176,9)) WHEN GTMED_S(176)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(177,9)) WHEN GTMED_S(177)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(178,9)) WHEN GTMED_S(178)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(179,9)) WHEN GTMED_S(179)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(180,9)) WHEN GTMED_S(180)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(181,9)) WHEN GTMED_S(181)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(182,9)) WHEN GTMED_S(182)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(183,9)) WHEN GTMED_S(183)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(184,9)) WHEN GTMED_S(184)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(185,9)) WHEN GTMED_S(185)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(186,9)) WHEN GTMED_S(186)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(187,9)) WHEN GTMED_S(187)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(188,9)) WHEN GTMED_S(188)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(189,9)) WHEN GTMED_S(189)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(190,9)) WHEN GTMED_S(190)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(191,9)) WHEN GTMED_S(191)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(192,9)) WHEN GTMED_S(192)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(193,9)) WHEN GTMED_S(193)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(194,9)) WHEN GTMED_S(194)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(195,9)) WHEN GTMED_S(195)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(196,9)) WHEN GTMED_S(196)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(197,9)) WHEN GTMED_S(197)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(198,9)) WHEN GTMED_S(198)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(199,9)) WHEN GTMED_S(199)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(200,9)) WHEN GTMED_S(200)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(201,9)) WHEN GTMED_S(201)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(202,9)) WHEN GTMED_S(202)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(203,9)) WHEN GTMED_S(203)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(204,9)) WHEN GTMED_S(204)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(205,9)) WHEN GTMED_S(205)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(206,9)) WHEN GTMED_S(206)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(207,9)) WHEN GTMED_S(207)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(208,9)) WHEN GTMED_S(208)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(209,9)) WHEN GTMED_S(209)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(210,9)) WHEN GTMED_S(210)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(211,9)) WHEN GTMED_S(211)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(212,9)) WHEN GTMED_S(212)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(213,9)) WHEN GTMED_S(213)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(214,9)) WHEN GTMED_S(214)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(215,9)) WHEN GTMED_S(215)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(216,9)) WHEN GTMED_S(216)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(217,9)) WHEN GTMED_S(217)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(218,9)) WHEN GTMED_S(218)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(219,9)) WHEN GTMED_S(219)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(220,9)) WHEN GTMED_S(220)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(221,9)) WHEN GTMED_S(221)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(222,9)) WHEN GTMED_S(222)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(223,9)) WHEN GTMED_S(223)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(224,9)) WHEN GTMED_S(224)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(225,9)) WHEN GTMED_S(225)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(226,9)) WHEN GTMED_S(226)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(227,9)) WHEN GTMED_S(227)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(228,9)) WHEN GTMED_S(228)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(229,9)) WHEN GTMED_S(229)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(230,9)) WHEN GTMED_S(230)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(231,9)) WHEN GTMED_S(231)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(232,9)) WHEN GTMED_S(232)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(233,9)) WHEN GTMED_S(233)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(234,9)) WHEN GTMED_S(234)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(235,9)) WHEN GTMED_S(235)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(236,9)) WHEN GTMED_S(236)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(237,9)) WHEN GTMED_S(237)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(238,9)) WHEN GTMED_S(238)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(239,9)) WHEN GTMED_S(239)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(240,9)) WHEN GTMED_S(240)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(241,9)) WHEN GTMED_S(241)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(242,9)) WHEN GTMED_S(242)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(243,9)) WHEN GTMED_S(243)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(244,9)) WHEN GTMED_S(244)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(245,9)) WHEN GTMED_S(245)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(246,9)) WHEN GTMED_S(246)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(247,9)) WHEN GTMED_S(247)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(248,9)) WHEN GTMED_S(248)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(249,9)) WHEN GTMED_S(249)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(250,9)) WHEN GTMED_S(250)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(251,9)) WHEN GTMED_S(251)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(252,9)) WHEN GTMED_S(252)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(253,9)) WHEN GTMED_S(253)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(254,9)) WHEN GTMED_S(254)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(255,9)) WHEN GTMED_S(255)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(256,9)) WHEN GTMED_S(256)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(257,9)) WHEN GTMED_S(257)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(258,9)) WHEN GTMED_S(258)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(259,9)) WHEN GTMED_S(259)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(260,9)) WHEN GTMED_S(260)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(261,9)) WHEN GTMED_S(261)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(262,9)) WHEN GTMED_S(262)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(263,9)) WHEN GTMED_S(263)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(264,9)) WHEN GTMED_S(264)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(265,9)) WHEN GTMED_S(265)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(266,9)) WHEN GTMED_S(266)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(267,9)) WHEN GTMED_S(267)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(268,9)) WHEN GTMED_S(268)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(269,9)) WHEN GTMED_S(269)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(270,9)) WHEN GTMED_S(270)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(271,9)) WHEN GTMED_S(271)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(272,9)) WHEN GTMED_S(272)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(273,9)) WHEN GTMED_S(273)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(274,9)) WHEN GTMED_S(274)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(275,9)) WHEN GTMED_S(275)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(276,9)) WHEN GTMED_S(276)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(277,9)) WHEN GTMED_S(277)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(278,9)) WHEN GTMED_S(278)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(279,9)) WHEN GTMED_S(279)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(280,9)) WHEN GTMED_S(280)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(281,9)) WHEN GTMED_S(281)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(282,9)) WHEN GTMED_S(282)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(283,9)) WHEN GTMED_S(283)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(284,9)) WHEN GTMED_S(284)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(285,9)) WHEN GTMED_S(285)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(286,9)) WHEN GTMED_S(286)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(287,9)) WHEN GTMED_S(287)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(288,9)) WHEN GTMED_S(288)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(289,9)) WHEN GTMED_S(289)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(290,9)) WHEN GTMED_S(290)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(291,9)) WHEN GTMED_S(291)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(292,9)) WHEN GTMED_S(292)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(293,9)) WHEN GTMED_S(293)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(294,9)) WHEN GTMED_S(294)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(295,9)) WHEN GTMED_S(295)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(296,9)) WHEN GTMED_S(296)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(297,9)) WHEN GTMED_S(297)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(298,9)) WHEN GTMED_S(298)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(299,9)) WHEN GTMED_S(299)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(300,9)) WHEN GTMED_S(300)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(301,9)) WHEN GTMED_S(301)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(302,9)) WHEN GTMED_S(302)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(303,9)) WHEN GTMED_S(303)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(304,9)) WHEN GTMED_S(304)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(305,9)) WHEN GTMED_S(305)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(306,9)) WHEN GTMED_S(306)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(307,9)) WHEN GTMED_S(307)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(308,9)) WHEN GTMED_S(308)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(309,9)) WHEN GTMED_S(309)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(310,9)) WHEN GTMED_S(310)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(311,9)) WHEN GTMED_S(311)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(312,9)) WHEN GTMED_S(312)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(313,9)) WHEN GTMED_S(313)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(314,9)) WHEN GTMED_S(314)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(315,9)) WHEN GTMED_S(315)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(316,9)) WHEN GTMED_S(316)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(317,9)) WHEN GTMED_S(317)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(318,9)) WHEN GTMED_S(318)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(319,9)) WHEN GTMED_S(319)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(320,9)) WHEN GTMED_S(320)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(321,9)) WHEN GTMED_S(321)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(322,9)) WHEN GTMED_S(322)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(323,9)) WHEN GTMED_S(323)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(324,9)) WHEN GTMED_S(324)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(325,9)) WHEN GTMED_S(325)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(326,9)) WHEN GTMED_S(326)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(327,9)) WHEN GTMED_S(327)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(328,9)) WHEN GTMED_S(328)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(329,9)) WHEN GTMED_S(329)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(330,9)) WHEN GTMED_S(330)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(331,9)) WHEN GTMED_S(331)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(332,9)) WHEN GTMED_S(332)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(333,9)) WHEN GTMED_S(333)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(334,9)) WHEN GTMED_S(334)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(335,9)) WHEN GTMED_S(335)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(336,9)) WHEN GTMED_S(336)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(337,9)) WHEN GTMED_S(337)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(338,9)) WHEN GTMED_S(338)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(339,9)) WHEN GTMED_S(339)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(340,9)) WHEN GTMED_S(340)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(341,9)) WHEN GTMED_S(341)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(342,9)) WHEN GTMED_S(342)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(343,9)) WHEN GTMED_S(343)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(344,9)) WHEN GTMED_S(344)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(345,9)) WHEN GTMED_S(345)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(346,9)) WHEN GTMED_S(346)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(347,9)) WHEN GTMED_S(347)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(348,9)) WHEN GTMED_S(348)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(349,9)) WHEN GTMED_S(349)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(350,9)) WHEN GTMED_S(350)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(351,9)) WHEN GTMED_S(351)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(352,9)) WHEN GTMED_S(352)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(353,9)) WHEN GTMED_S(353)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(354,9)) WHEN GTMED_S(354)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(355,9)) WHEN GTMED_S(355)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(356,9)) WHEN GTMED_S(356)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(357,9)) WHEN GTMED_S(357)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(358,9)) WHEN GTMED_S(358)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(359,9)) WHEN GTMED_S(359)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(360,9)) WHEN GTMED_S(360)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(361,9)) WHEN GTMED_S(361)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(362,9)) WHEN GTMED_S(362)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(363,9)) WHEN GTMED_S(363)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(364,9)) WHEN GTMED_S(364)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(365,9)) WHEN GTMED_S(365)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(366,9)) WHEN GTMED_S(366)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(367,9)) WHEN GTMED_S(367)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(368,9)) WHEN GTMED_S(368)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(369,9)) WHEN GTMED_S(369)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(370,9)) WHEN GTMED_S(370)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(371,9)) WHEN GTMED_S(371)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(372,9)) WHEN GTMED_S(372)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(373,9)) WHEN GTMED_S(373)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(374,9)) WHEN GTMED_S(374)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(375,9)) WHEN GTMED_S(375)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(376,9)) WHEN GTMED_S(376)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(377,9)) WHEN GTMED_S(377)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(378,9)) WHEN GTMED_S(378)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(379,9)) WHEN GTMED_S(379)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(380,9)) WHEN GTMED_S(380)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(381,9)) WHEN GTMED_S(381)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(382,9)) WHEN GTMED_S(382)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(383,9)) WHEN GTMED_S(383)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(384,9)) WHEN GTMED_S(384)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(385,9)) WHEN GTMED_S(385)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(386,9)) WHEN GTMED_S(386)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(387,9)) WHEN GTMED_S(387)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(388,9)) WHEN GTMED_S(388)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(389,9)) WHEN GTMED_S(389)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(390,9)) WHEN GTMED_S(390)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(391,9)) WHEN GTMED_S(391)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(392,9)) WHEN GTMED_S(392)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(393,9)) WHEN GTMED_S(393)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(394,9)) WHEN GTMED_S(394)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(395,9)) WHEN GTMED_S(395)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(396,9)) WHEN GTMED_S(396)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(397,9)) WHEN GTMED_S(397)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(398,9)) WHEN GTMED_S(398)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(399,9)) WHEN GTMED_S(399)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(400,9)) WHEN GTMED_S(400)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(401,9)) WHEN GTMED_S(401)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(402,9)) WHEN GTMED_S(402)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(403,9)) WHEN GTMED_S(403)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(404,9)) WHEN GTMED_S(404)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(405,9)) WHEN GTMED_S(405)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(406,9)) WHEN GTMED_S(406)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(407,9)) WHEN GTMED_S(407)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(408,9)) WHEN GTMED_S(408)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(409,9)) WHEN GTMED_S(409)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(410,9)) WHEN GTMED_S(410)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(411,9)) WHEN GTMED_S(411)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(412,9)) WHEN GTMED_S(412)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(413,9)) WHEN GTMED_S(413)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(414,9)) WHEN GTMED_S(414)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(415,9)) WHEN GTMED_S(415)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(416,9)) WHEN GTMED_S(416)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(417,9)) WHEN GTMED_S(417)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(418,9)) WHEN GTMED_S(418)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(419,9)) WHEN GTMED_S(419)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(420,9)) WHEN GTMED_S(420)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(421,9)) WHEN GTMED_S(421)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(422,9)) WHEN GTMED_S(422)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(423,9)) WHEN GTMED_S(423)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(424,9)) WHEN GTMED_S(424)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(425,9)) WHEN GTMED_S(425)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(426,9)) WHEN GTMED_S(426)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(427,9)) WHEN GTMED_S(427)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(428,9)) WHEN GTMED_S(428)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(429,9)) WHEN GTMED_S(429)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(430,9)) WHEN GTMED_S(430)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(431,9)) WHEN GTMED_S(431)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(432,9)) WHEN GTMED_S(432)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(433,9)) WHEN GTMED_S(433)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(434,9)) WHEN GTMED_S(434)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(435,9)) WHEN GTMED_S(435)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(436,9)) WHEN GTMED_S(436)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(437,9)) WHEN GTMED_S(437)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(438,9)) WHEN GTMED_S(438)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(439,9)) WHEN GTMED_S(439)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(440,9)) WHEN GTMED_S(440)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(441,9)) WHEN GTMED_S(441)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(442,9)) WHEN GTMED_S(442)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(443,9)) WHEN GTMED_S(443)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(444,9)) WHEN GTMED_S(444)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(445,9)) WHEN GTMED_S(445)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(446,9)) WHEN GTMED_S(446)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(447,9)) WHEN GTMED_S(447)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(448,9)) WHEN GTMED_S(448)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(449,9)) WHEN GTMED_S(449)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(450,9)) WHEN GTMED_S(450)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(451,9)) WHEN GTMED_S(451)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(452,9)) WHEN GTMED_S(452)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(453,9)) WHEN GTMED_S(453)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(454,9)) WHEN GTMED_S(454)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(455,9)) WHEN GTMED_S(455)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(456,9)) WHEN GTMED_S(456)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(457,9)) WHEN GTMED_S(457)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(458,9)) WHEN GTMED_S(458)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(459,9)) WHEN GTMED_S(459)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(460,9)) WHEN GTMED_S(460)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(461,9)) WHEN GTMED_S(461)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(462,9)) WHEN GTMED_S(462)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(463,9)) WHEN GTMED_S(463)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(464,9)) WHEN GTMED_S(464)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(465,9)) WHEN GTMED_S(465)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(466,9)) WHEN GTMED_S(466)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(467,9)) WHEN GTMED_S(467)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(468,9)) WHEN GTMED_S(468)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(469,9)) WHEN GTMED_S(469)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(470,9)) WHEN GTMED_S(470)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(471,9)) WHEN GTMED_S(471)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(472,9)) WHEN GTMED_S(472)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(473,9)) WHEN GTMED_S(473)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(474,9)) WHEN GTMED_S(474)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(475,9)) WHEN GTMED_S(475)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(476,9)) WHEN GTMED_S(476)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(477,9)) WHEN GTMED_S(477)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(478,9)) WHEN GTMED_S(478)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(479,9)) WHEN GTMED_S(479)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(480,9)) WHEN GTMED_S(480)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(481,9)) WHEN GTMED_S(481)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(482,9)) WHEN GTMED_S(482)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(483,9)) WHEN GTMED_S(483)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(484,9)) WHEN GTMED_S(484)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(485,9)) WHEN GTMED_S(485)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(486,9)) WHEN GTMED_S(486)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(487,9)) WHEN GTMED_S(487)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(488,9)) WHEN GTMED_S(488)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(489,9)) WHEN GTMED_S(489)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(490,9)) WHEN GTMED_S(490)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(491,9)) WHEN GTMED_S(491)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(492,9)) WHEN GTMED_S(492)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(493,9)) WHEN GTMED_S(493)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(494,9)) WHEN GTMED_S(494)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(495,9)) WHEN GTMED_S(495)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(496,9)) WHEN GTMED_S(496)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(497,9)) WHEN GTMED_S(497)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(498,9)) WHEN GTMED_S(498)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(499,9)) WHEN GTMED_S(499)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(500,9)) WHEN GTMED_S(500)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(501,9)) WHEN GTMED_S(501)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(502,9)) WHEN GTMED_S(502)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(503,9)) WHEN GTMED_S(503)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(504,9)) WHEN GTMED_S(504)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(505,9)) WHEN GTMED_S(505)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(506,9)) WHEN GTMED_S(506)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(507,9)) WHEN GTMED_S(507)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(508,9)) WHEN GTMED_S(508)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(509,9)) WHEN GTMED_S(509)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(510,9)) WHEN GTMED_S(510)='1' ELSE
				 STD_LOGIC_VECTOR(TO_UNSIGNED(511,9)) WHEN GTMED_S(511)='1' ELSE (OTHERS=>'0');
				 
				 

END ARCHITECTURE RTL;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

--9 BIT DECODER
ENTITY SELECTORBIN IS 
PORT( SEL: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		ENABLE: IN STD_LOGIC;
		LUT_OUT: OUT STD_LOGIC_VECTOR (511 DOWNTO 0)
		);
END ENTITY SELECTORBIN;

ARCHITECTURE RTL OF SELECTORBIN IS
BEGIN
DECO:PROCESS(SEL,ENABLE)
BEGIN
IF(ENABLE='0') THEN 
CASE TO_INTEGER(UNSIGNED(SEL)) IS
WHEN 0 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
WHEN 1 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";
WHEN 2 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC";
WHEN 3 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8";
WHEN 4 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0";
WHEN 5 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0";
WHEN 6 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0";
WHEN 7 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80";
WHEN 8 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00";
WHEN 9 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00";
WHEN 10 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00";
WHEN 11 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800";
WHEN 12 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000";
WHEN 13 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000";
WHEN 14 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000";
WHEN 15 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000";
WHEN 16 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000";
WHEN 17 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000";
WHEN 18 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000";
WHEN 19 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000";
WHEN 20 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000";
WHEN 21 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000";
WHEN 22 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000";
WHEN 23 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000";
WHEN 24 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000";
WHEN 25 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000";
WHEN 26 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000";
WHEN 27 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000";
WHEN 28 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000";
WHEN 29 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000";
WHEN 30 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000";
WHEN 31 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000";
WHEN 32 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000";
WHEN 33 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000";
WHEN 34 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000";
WHEN 35 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000";
WHEN 36 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000";
WHEN 37 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000";
WHEN 38 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000";
WHEN 39 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000";
WHEN 40 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000";
WHEN 41 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000";
WHEN 42 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000";
WHEN 43 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000";
WHEN 44 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000";
WHEN 45 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000";
WHEN 46 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000";
WHEN 47 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000";
WHEN 48 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000";
WHEN 49 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000";
WHEN 50 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000";
WHEN 51 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000";
WHEN 52 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000";
WHEN 53 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000";
WHEN 54 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000";
WHEN 55 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000";
WHEN 56 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000";
WHEN 57 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000";
WHEN 58 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000";
WHEN 59 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000";
WHEN 60 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000";
WHEN 61 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000";
WHEN 62 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000";
WHEN 63 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000";
WHEN 64 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000";
WHEN 65 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000";
WHEN 66 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000";
WHEN 67 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000";
WHEN 68 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000";
WHEN 69 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000";
WHEN 70 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000";
WHEN 71 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000";
WHEN 72 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000";
WHEN 73 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000";
WHEN 74 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000";
WHEN 75 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000";
WHEN 76 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000";
WHEN 77 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000";
WHEN 78 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000";
WHEN 79 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000";
WHEN 80 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000";
WHEN 81 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
WHEN 82 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000";
WHEN 83 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000";
WHEN 84 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000";
WHEN 85 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000";
WHEN 86 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000";
WHEN 87 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
WHEN 88 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
WHEN 89 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000";
WHEN 90 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000";
WHEN 91 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000";
WHEN 92 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000";
WHEN 93 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000";
WHEN 94 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000";
WHEN 95 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000";
WHEN 96 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000";
WHEN 97 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000";
WHEN 98 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000";
WHEN 99 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000";
WHEN 100 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000";
WHEN 101 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000";
WHEN 102 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000";
WHEN 103 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000";
WHEN 104 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000";
WHEN 105 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000";
WHEN 106 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000";
WHEN 107 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000";
WHEN 108 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000";
WHEN 109 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000";
WHEN 110 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000";
WHEN 111 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000";
WHEN 112 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000";
WHEN 113 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000";
WHEN 114 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000";
WHEN 115 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000";
WHEN 116 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000";
WHEN 117 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000";
WHEN 118 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000";
WHEN 119 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000";
WHEN 120 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000";
WHEN 121 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000";
WHEN 122 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000";
WHEN 123 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000";
WHEN 124 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000";
WHEN 125 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000";
WHEN 126 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000";
WHEN 127 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000";
WHEN 128 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000";
WHEN 129 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000";
WHEN 130 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000";
WHEN 131 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000";
WHEN 132 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000";
WHEN 133 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000";
WHEN 134 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000";
WHEN 135 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000";
WHEN 136 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000";
WHEN 137 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000";
WHEN 138 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000";
WHEN 139 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000";
WHEN 140 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000";
WHEN 141 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000";
WHEN 142 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000";
WHEN 143 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000";
WHEN 144 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000";
WHEN 145 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000";
WHEN 146 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000";
WHEN 147 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000";
WHEN 148 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000";
WHEN 149 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000";
WHEN 150 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000";
WHEN 151 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000";
WHEN 152 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000";
WHEN 153 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000";
WHEN 154 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000";
WHEN 155 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000";
WHEN 156 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000";
WHEN 157 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000";
WHEN 158 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000";
WHEN 159 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000";
WHEN 160 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000";
WHEN 161 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000";
WHEN 162 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000";
WHEN 163 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000";
WHEN 164 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000";
WHEN 165 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000";
WHEN 166 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000";
WHEN 167 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000";
WHEN 168 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000";
WHEN 169 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000";
WHEN 170 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000";
WHEN 171 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000";
WHEN 172 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000";
WHEN 173 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000";
WHEN 174 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000";
WHEN 175 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000";
WHEN 176 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000";
WHEN 177 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000";
WHEN 178 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000";
WHEN 179 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000";
WHEN 180 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000";
WHEN 181 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000";
WHEN 182 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000";
WHEN 183 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000";
WHEN 184 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000";
WHEN 185 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000";
WHEN 186 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000";
WHEN 187 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000";
WHEN 188 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000";
WHEN 189 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000";
WHEN 190 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000";
WHEN 191 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000";
WHEN 192 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000";
WHEN 193 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000";
WHEN 194 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000";
WHEN 195 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000";
WHEN 196 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000";
WHEN 197 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000";
WHEN 198 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000";
WHEN 199 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000";
WHEN 200 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000";
WHEN 201 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000";
WHEN 202 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000";
WHEN 203 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000";
WHEN 204 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000";
WHEN 205 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000";
WHEN 206 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000";
WHEN 207 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000";
WHEN 208 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000";
WHEN 209 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000";
WHEN 210 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000";
WHEN 211 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000";
WHEN 212 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000";
WHEN 213 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000";
WHEN 214 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000";
WHEN 215 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000";
WHEN 216 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000";
WHEN 217 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000";
WHEN 218 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000";
WHEN 219 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000";
WHEN 220 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000";
WHEN 221 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000";
WHEN 222 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000";
WHEN 223 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000";
WHEN 224 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000";
WHEN 225 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000";
WHEN 226 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000";
WHEN 227 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000";
WHEN 228 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000";
WHEN 229 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000";
WHEN 230 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000";
WHEN 231 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000";
WHEN 232 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000";
WHEN 233 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000";
WHEN 234 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000";
WHEN 235 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000";
WHEN 236 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000";
WHEN 237 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000";
WHEN 238 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000";
WHEN 239 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000";
WHEN 240 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000";
WHEN 241 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000";
WHEN 242 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000";
WHEN 243 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000";
WHEN 244 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000";
WHEN 245 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000";
WHEN 246 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000";
WHEN 247 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000";
WHEN 248 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000";
WHEN 249 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000";
WHEN 250 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000";
WHEN 251 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000";
WHEN 252 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000";
WHEN 253 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000";
WHEN 254 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000";
WHEN 255 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000";
WHEN 256 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000";
WHEN 257 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000";
WHEN 258 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000";
WHEN 259 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000";
WHEN 260 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000";
WHEN 261 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000";
WHEN 262 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000";
WHEN 263 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000";
WHEN 264 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000";
WHEN 265 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000";
WHEN 266 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000";
WHEN 267 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000";
WHEN 268 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000";
WHEN 269 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000";
WHEN 270 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000";
WHEN 271 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000";
WHEN 272 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000";
WHEN 273 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000";
WHEN 274 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000";
WHEN 275 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000";
WHEN 276 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 277 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 278 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 279 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 280 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 281 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 282 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 283 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 284 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 285 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 286 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 287 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 288 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 289 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 290 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 291 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 292 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 293 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 294 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 295 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 296 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 297 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 298 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 299 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 300 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 301 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 302 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 303 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 304 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 305 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 306 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 307 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 308 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 309 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 310 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 311 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 312 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 313 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 314 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 315 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 316 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 317 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 318 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 319 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 320 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 321 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 322 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 323 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 324 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 325 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 326 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 327 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 328 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 329 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 330 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 331 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 332 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 333 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 334 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 335 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 336 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 337 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 338 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 339 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 340 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 341 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 342 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 343 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 344 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 345 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 346 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 347 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 348 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 349 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 350 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 351 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 352 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 353 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 354 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 355 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 356 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 357 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 358 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 359 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 360 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 361 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 362 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 363 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 364 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 365 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 366 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 367 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 368 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 369 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 370 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 371 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 372 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 373 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 374 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 375 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 376 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 377 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 378 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 379 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 380 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 381 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 382 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 383 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 384 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 385 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 386 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 387 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 388 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 389 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 390 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 391 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 392 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 393 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 394 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 395 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 396 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 397 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 398 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 399 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 400 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 401 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 402 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 403 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 404 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 405 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 406 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 407 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 408 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 409 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 410 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 411 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 412 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 413 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 414 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 415 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 416 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 417 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 418 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 419 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 420 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 421 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 422 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 423 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 424 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 425 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 426 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 427 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 428 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 429 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 430 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 431 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 432 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 433 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 434 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 435 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 436 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 437 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 438 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 439 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 440 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 441 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 442 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 443 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 444 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 445 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 446 =>LUT_OUT<= X"FFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 447 =>LUT_OUT<= X"FFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 448 =>LUT_OUT<= X"FFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 449 =>LUT_OUT<= X"FFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 450 =>LUT_OUT<= X"FFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 451 =>LUT_OUT<= X"FFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 452 =>LUT_OUT<= X"FFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 453 =>LUT_OUT<= X"FFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 454 =>LUT_OUT<= X"FFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 455 =>LUT_OUT<= X"FFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 456 =>LUT_OUT<= X"FFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 457 =>LUT_OUT<= X"FFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 458 =>LUT_OUT<= X"FFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 459 =>LUT_OUT<= X"FFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 460 =>LUT_OUT<= X"FFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 461 =>LUT_OUT<= X"FFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 462 =>LUT_OUT<= X"FFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 463 =>LUT_OUT<= X"FFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 464 =>LUT_OUT<= X"FFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 465 =>LUT_OUT<= X"FFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 466 =>LUT_OUT<= X"FFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 467 =>LUT_OUT<= X"FFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 468 =>LUT_OUT<= X"FFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 469 =>LUT_OUT<= X"FFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 470 =>LUT_OUT<= X"FFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 471 =>LUT_OUT<= X"FFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 472 =>LUT_OUT<= X"FFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 473 =>LUT_OUT<= X"FFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 474 =>LUT_OUT<= X"FFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 475 =>LUT_OUT<= X"FFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 476 =>LUT_OUT<= X"FFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 477 =>LUT_OUT<= X"FFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 478 =>LUT_OUT<= X"FFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 479 =>LUT_OUT<= X"FFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 480 =>LUT_OUT<= X"FFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 481 =>LUT_OUT<= X"FFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 482 =>LUT_OUT<= X"FFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 483 =>LUT_OUT<= X"FFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 484 =>LUT_OUT<= X"FFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 485 =>LUT_OUT<= X"FFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 486 =>LUT_OUT<= X"FFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 487 =>LUT_OUT<= X"FFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 488 =>LUT_OUT<= X"FFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 489 =>LUT_OUT<= X"FFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 490 =>LUT_OUT<= X"FFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 491 =>LUT_OUT<= X"FFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 492 =>LUT_OUT<= X"FFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 493 =>LUT_OUT<= X"FFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 494 =>LUT_OUT<= X"FFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 495 =>LUT_OUT<= X"FFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 496 =>LUT_OUT<= X"FFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 497 =>LUT_OUT<= X"FFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 498 =>LUT_OUT<= X"FFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 499 =>LUT_OUT<= X"FFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 500 =>LUT_OUT<= X"FFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 501 =>LUT_OUT<= X"FFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 502 =>LUT_OUT<= X"FFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 503 =>LUT_OUT<= X"FF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 504 =>LUT_OUT<= X"FF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 505 =>LUT_OUT<= X"FE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 506 =>LUT_OUT<= X"FC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 507 =>LUT_OUT<= X"F8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 508 =>LUT_OUT<= X"F0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 509 =>LUT_OUT<= X"E0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 510 =>LUT_OUT<= X"C0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN 511 =>LUT_OUT<= X"80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
WHEN OTHERS =>LUT_OUT<= (OTHERS=>'0');
END CASE;
ELSE
LUT_OUT<=(OTHERS=>'0');
END IF;

END PROCESS DECO;
END ARCHITECTURE RTL;
